`timescale 1ns / 1ps

module receiver #(
    parameter CLKS_PER_BIT = 217
)(
    input  wire        			CLK,
    input  wire        			Rx_in,
    output wire        			Rx_DV_out,
    output wire [7:0]  			Rx_Byte_out
);

    //==================================================//
    //                 State Encoding                   //
    //==================================================//
    localparam s_IDLE         	= 3'b000;
    localparam s_RX_START_BIT 	= 3'b001;
    localparam s_RX_DATA_BITS 	= 3'b010;
    localparam s_RX_STOP_BIT  	= 3'b011;
    localparam s_CLEANUP      	= 3'b100;

    //==================================================//
    //                   Registers                      //
    //==================================================//
    reg           Rx_Data_R_r   = 1'b1;
    reg           Rx_Data_r     = 1'b1;
    reg  [7:0]    Clock_Count_r = 0;
    reg  [2:0]    Bit_Index_r   = 0;
    reg  [7:0]    Rx_Byte_r     = 0;
    reg           Rx_DV_r       = 0;
	
	reg  [7:0]    LED_r			= 0;

    reg  [2:0]    current_state_r = s_IDLE;   // current state
    reg  [2:0]    next_state_r;    // next state

    //==================================================//
    //             Input Synchronization                //
    //==================================================//
    always @(posedge CLK) begin
        Rx_Data_R_r <= Rx_in;
        Rx_Data_r   <= Rx_Data_R_r;
    end

    //==================================================//
    //                  Next State Logic                //
    //==================================================//
    always @* begin
        case (current_state_r)
            s_IDLE:
                if (Rx_Data_r == 1'b0)
                    next_state_r = s_RX_START_BIT;
                else
                    next_state_r = s_IDLE;

            s_RX_START_BIT:
                if (Clock_Count_r == (CLKS_PER_BIT - 1) / 2)
                    if (Rx_Data_r == 1'b0)
                        next_state_r = s_RX_DATA_BITS;
                    else
                        next_state_r = s_IDLE;
                else
                    next_state_r = s_RX_START_BIT;

            s_RX_DATA_BITS:
                if (Clock_Count_r < CLKS_PER_BIT - 1)
                    next_state_r = s_RX_DATA_BITS;
                else if (Bit_Index_r < 7)
                    next_state_r = s_RX_DATA_BITS;
                else
                    next_state_r = s_RX_STOP_BIT;

            s_RX_STOP_BIT:
                if (Clock_Count_r < CLKS_PER_BIT - 1)
                    next_state_r = s_RX_STOP_BIT;
                else
                    next_state_r = s_CLEANUP;

            s_CLEANUP:
                next_state_r = s_IDLE;

            default:
                next_state_r = s_IDLE;
        endcase
    end

    //==================================================//
    //                State Register (FSM)              //
    //==================================================//
    always @(posedge CLK) begin
        current_state_r <= next_state_r;
    end

    //==================================================//
    //                   Datapath                       //
    //==================================================//
    always @(posedge CLK) begin
        case (current_state_r)
            s_IDLE: begin
                Rx_DV_r       <= 1'b0;
                Clock_Count_r <= 0;
                Bit_Index_r   <= 0;
            end

            s_RX_START_BIT: begin
                if (Clock_Count_r == (CLKS_PER_BIT - 1) / 2) begin
                    if (Rx_Data_r == 1'b0)
                        Clock_Count_r <= 0;
                end else
                    Clock_Count_r <= Clock_Count_r + 1;
            end

            s_RX_DATA_BITS: begin
                if (Clock_Count_r < CLKS_PER_BIT - 1) begin
                    Clock_Count_r <= Clock_Count_r + 1;
                end else begin
                    Clock_Count_r          <= 0;
                    Rx_Byte_r[Bit_Index_r] <= Rx_Data_r;
                    if (Bit_Index_r < 7)
                        Bit_Index_r <= Bit_Index_r + 1;
                    else
                        Bit_Index_r <= 0;
                end
            end

            s_RX_STOP_BIT: begin
                if (Clock_Count_r < CLKS_PER_BIT - 1) begin
                    Clock_Count_r <= Clock_Count_r + 1;
                end else begin
                    Rx_DV_r       <= 1'b1;
                    Clock_Count_r <= 0;
                end
            end

            s_CLEANUP: begin
                Rx_DV_r <= 1'b0;
            end

            default: begin
                Rx_DV_r       <= 1'b0;
                Clock_Count_r <= 0;
                Bit_Index_r   <= 0;
            end
        endcase
    end

    //==================================================//
    //                     Output                       //
    //==================================================//
    assign Rx_DV_out   = Rx_DV_r;
    assign Rx_Byte_out = Rx_Byte_r;

endmodule
