// add_tb_pkg.sv
package add_tb_pkg;
    `include "packet.sv"
    `include "Simulus.sv"
    `include "Driver.sv"
    `include "Monitor.sv"
    `include "Scoreboard.sv"
endpackage
